LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CLK_ABAJO is
    Port ( CLK : in  STD_LOGIC;
           CLKOUT : out  STD_LOGIC);
end CLK_ABAJO;

architecture Behavioral of CLK_ABAJO is
	SIGNAL CLK25: STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL SALIDA : STD_LOGIC;
begin
	-- RELOJ DE 25MHZ
	PROCESS (CLK)
		BEGIN
		IF CLK'EVENT AND CLK='1' THEN
			IF CLK25 = "1000" THEN
				CLK25 <= "0000";
				SALIDA <= NOT SALIDA;
			ELSE
				CLK25 <= CLK25 + 1;
		ELSE NULL;
		END IF;
	END PROCESS;
	
	CLKOUT <= SALIDA;

end Behavioral;

