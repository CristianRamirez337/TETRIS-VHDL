LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEBOUNCE IS
	PORT (
		CLK : IN STD_LOGIC;
		DIN : IN STD_LOGIC;
		QOUT : OUT STD_LOGIC);
END DEBOUNCE;

ARCHITECTURE Behavioral OF DEBOUNCE IS
	SIGNAL Q1, Q2, Q3 : STD_LOGIC;
BEGIN
	PROCESS (CLK)
	BEGIN
		IF (CLK = '1' AND CLK'EVENT) THEN
			Q1 <= DIN;
			Q2 <= Q1;
			Q3 <= Q2;
		END IF;
	END PROCESS;

	QOUT <= Q1 AND Q2 AND NOT Q3;

END Behavioral;