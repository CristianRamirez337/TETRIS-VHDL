LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CLK_500HZ IS
	PORT (
		MCLK : IN STD_LOGIC;
		CLKOUT : OUT STD_LOGIC
	);
END CLK_500HZ;

ARCHITECTURE Behavioral OF CLK_500HZ IS
	SIGNAL COUNTER : INTEGER RANGE 0 TO 49_999 := 0;
	SIGNAL C500HZ : STD_LOGIC;
BEGIN
	PROCESS (MCLK)
	BEGIN
		IF MCLK = '1' AND MCLK'EVENT THEN
			IF COUNTER = 49_999 THEN
				COUNTER <= 0;
				C500HZ <= NOT C500HZ;
			ELSE COUNTER <= COUNTER + 1;
			END IF;
		ELSE NULL;
		END IF;
	END PROCESS;

	CLKOUT <= C500HZ;
END Behavioral;