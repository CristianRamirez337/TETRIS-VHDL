LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECODER IS
	PORT(
		HS,VS: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		HS_OUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		VS_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END DECODER;

ARCHITECTURE Behavioral OF DECODER IS

BEGIN
	PROCESS(HS) --X(150,640), Y(50,480) 
		BEGIN
			IF (HS > "0100101100" and HS <  "0100111011") THEN
				HS_OUT <= "0001";
			ELSIF (HS > "0100111011" and HS <  "0101001010") THEN
				HS_OUT <= "0010";
			ELSIF (HS > "0101001010" and HS <  "0101011001") THEN
				HS_OUT <= "0011";
			ELSIF (HS > "0101011001" and HS <  "0101101000") THEN
				HS_OUT <= "0100";
			ELSIF (HS > "0101101000" and HS <  "0101110111") THEN
				HS_OUT <= "0101";
			ELSIF (HS > "0101110111" and HS <  "0110000110") THEN
				HS_OUT <= "0110";
			ELSIF (HS > "0110000110" and HS <  "0110010101") THEN
				HS_OUT <= "0111";
			ELSIF (HS > "0110010101" and HS <  "0110100100") THEN
				HS_OUT <= "1000";
			ELSIF (HS > "0110100100" and HS <  "0110110011") THEN
				HS_OUT <= "1001";
			ELSIF (HS > "0110110011" and HS <  "0111000010") THEN
				HS_OUT <= "1010";
			ELSE
				HS_OUT <= "0000";
			END IF;
	END PROCESS;
	
	PROCESS(VS) --X(150,640), Y(50,480) 
		BEGIN
			IF (VS > "0011000011" and VS <  "0011010010") THEN
				VS_OUT <= "00001";
			ELSIF (VS > "0011010010" and VS <  "0011100001") THEN
				VS_OUT <= "00010";
			ELSIF (VS > "0011100001" and VS <  "0011110000") THEN
				VS_OUT <= "00011";
			ELSIF (VS > "0011110000" and VS <  "0011111111") THEN
				VS_OUT <= "00100";
			ELSIF (VS > "0011111111" and VS <  "0100001110") THEN -- Vertical 0,1
				VS_OUT <= "00101";
			ELSIF (VS > "0100001110" and VS <  "0100011101") THEN
				VS_OUT <= "00110";
			ELSIF (VS > "0100011101" and VS <  "0100101100") THEN
				VS_OUT <= "00111";
			ELSIF (VS > "0100101100" and VS <  "0100111011") THEN
				VS_OUT <= "01000";
			ELSIF (VS > "0100111011" and VS <  "0101001010") THEN
				VS_OUT <= "01001";
			ELSIF (VS > "0101001010" and VS <  "0101011001") THEN
				VS_OUT <= "01010";
			ELSIF (VS > "0101011001" and VS <  "0101101000") THEN
				VS_OUT <= "01011";
			ELSIF (VS > "0101101000" and VS <  "0101110111") THEN
				VS_OUT <= "01100";
			ELSIF (VS > "0101110111" and VS <  "0110000110") THEN
				VS_OUT <= "01101";
			ELSIF (VS > "0110000110" and VS <  "0110010101") THEN
				VS_OUT <= "01110";
			ELSIF (VS > "0110010101" and VS <  "0110100100") THEN
				VS_OUT <= "01111";
			ELSIF (VS > "0110100100" and VS <  "0110110011") THEN -- Desde aqui correcciones lado derecho
				VS_OUT <= "10000";
			ELSIF (VS > "0110110011" and VS <  "0111000010") THEN
				VS_OUT <= "10001";
			ELSIF (VS > "0111000010" and VS <  "0111010001") THEN
				VS_OUT <= "10010";
			ELSIF (VS > "0111010001" and VS <  "0111100000") THEN
				VS_OUT <= "10011";
			ELSE
				VS_OUT <= "00000";
			END IF;
	END PROCESS;
END Behavioral;